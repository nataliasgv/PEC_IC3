library IEEE;
use IEEE.std_logic_1164.all;


-- esta entity sirve para la architecture ej1a y ej1b
entity ej1 is
port( F, G : out std_logic;
x, y, z : in std_logic);
end entity ej1;


