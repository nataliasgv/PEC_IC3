library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
	
entity AND_gate is
	port (
		A, B : in std_logic;
		Y : out std_logic
	);
end entity AND_gate;
	
architecture estructuraAND of AND_gate is
begin
	Y <= A and B;
end architecture estructuraAND;
